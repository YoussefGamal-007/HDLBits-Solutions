module top_module (
    output out);

    supply0 GND;
    assign out = GND;
endmodule
