module top_module( output one );

// Insert your code here
    supply1 VDD;
    assign one = VDD ;

endmodule
